module MUL(a, b)