module Xor_1(a,b,y);
input logic a, b;
output logic y;
assign y = a^b;
endmodule
